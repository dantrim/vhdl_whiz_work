entity T06_SignalTb is
end entity;

architecture sim of T06_SignalTb is

    -- TODO: Declare a signal of type integer with initial value 0

begin

    process is
        -- TODO: Declare a variable of type integer with initial value 0
    begin

        report "*** Process begin ***";

        -- TODO: Increment the signal and variable here

        -- TODO: Print the signal and variable values here

        -- TODO: Increment the signal and variable here

        -- TODO: Print the signal and variable values here

        wait for 10 ns;

        -- TODO: Print the signal and variable values here

    end process;

end architecture;