library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- TODO: Create an entity with a port declaration
--       
--       The entity name shall be T15_Mux
--
--       The port shall have 5 inputs of type unsigned:
--       Sig1, Sig2, Sig3, Sig4, and Sel
--       And one output of type unsigned: Output

architecture rtl of T15_Mux is
begin

    -- TODO: Move the MUX process from T15_PortMap.vhd to here
    
end architecture;