library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity T17_FlipFlop is
port(
    -- TODO: Complete the port of a flip flop.
    --       
    --       The inputs of type std_logic shall be:
    --          Clk (clock)
    --          nRst (negative reset)
    --          Input
    --
    --       The output of type std_logic shall be: Output
);
end entity;

architecture rtl of T17_FlipFlop is
begin

    -- Flip-flop with synchronized reset
    -- TODO: Implement a Flip-flop in a clocked process here.
    --       Use negative synchronous reset.

end architecture;