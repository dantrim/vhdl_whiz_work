entity T04_ForLoopTb is
end entity;

architecture sim of T04_ForLoopTb is
begin

    process is
    begin

        -- TASK: Create For-loop here.
        --       Print the value of the implicit variable inside of the loop
        
        wait;

    end process;

end architecture;